// Copyright 2021 ETH Zurich and University of Bologna.
// Solderpad Hardware License, Version 0.51, see LICENSE for details.
// SPDX-License-Identifier: SHL-0.51
//
// Author: Matheus Cavalcante <matheusd@iis.ee.ethz.ch>
// Description:
// This is the vector register file of one lane.

module vector_regfile import ara_pkg::*; #(
    parameter  int  unsigned NrBanks   = 0,     // Number of banks in the vector register file
    parameter  int  unsigned VRFSize   = 0,     // Size of the VRF, in bits
    parameter  type          vaddr_t   = logic,
    // Dependant parameters. DO NOT CHANGE!
    localparam int  unsigned DataWidth = $bits(elen_t),
    localparam int  unsigned StrbWidth = DataWidth / 8,
    localparam type          strb_t    = logic [StrbWidth-1:0]
  ) (
    input  logic                           clk_i,
    input  logic                           rst_ni,
    // Interface with the VRF
    input  logic     [NrBanks-1:0]         req_i,
    input  vaddr_t   [NrBanks-1:0]         addr_i,
    input  opqueue_e [NrBanks-1:0]         tgt_opqueue_i,
    input  logic     [NrBanks-1:0]         wen_i,
    input  elen_t    [NrBanks-1:0]         wdata_i,
    input  strb_t    [NrBanks-1:0]         be_i,
    // Operands
    output elen_t    [NrOperandQueues-1:0] operand_o,
    output logic     [NrOperandQueues-1:0] operand_valid_o
  );

`include "common_cells/registers.svh"

  //////////////////
  //  Parameters  //
  //////////////////

  localparam int unsigned NumWords = VRFSize / NrBanks / DataWidth;

  ///////////////
  //  Signals  //
  ///////////////

  elen_t    [NrBanks-1:0] rdata;
  logic     [NrBanks-1:0] rdata_valid_q;
  opqueue_e [NrBanks-1:0] tgt_opqueue_q;

  // Generate the rdata_valid and tgt_opqueue signals by delaying the request by one cycle
  always_ff @(posedge clk_i or negedge rst_ni) begin: p_rdata_valid
    if (!rst_ni) begin
      rdata_valid_q <= '0;
      tgt_opqueue_q <= '0;
    end else begin
      rdata_valid_q <= req_i & ~wen_i;
      tgt_opqueue_q <= tgt_opqueue_i;
    end
  end

  /////////////
  //  Banks  //
  /////////////

  for (genvar bank = 0; bank < NrBanks; bank++) begin: gen_banks
`ifndef VERILATOR
    // Clock gate
    logic vrf_clk;
    logic sram_active_q;
    `FF(sram_active_q, req_i[bank], 1'b0)

    tc_clk_gating i_vrf_ckg (
      .clk_i    (clk_i                       ),
      .test_en_i(1'b0                        ),
      .en_i     (req_i[bank] || sram_active_q),
      .clk_o    (vrf_clk                     )
    );
`else
    logic vrf_clk;

    assign vrf_clk = clk_i;
`endif

`ifndef TARGET_SRAM_MC
    tc_sram #(
      .NumWords (NumWords ),
      .DataWidth(DataWidth),
      .NumPorts (1        )
    ) data_sram (
      .clk_i  (vrf_clk                           ),
      .rst_ni (rst_ni                            ),
      .req_i  (req_i[bank]                       ),
      .we_i   (wen_i[bank]                       ),
      .rdata_o(rdata[bank]                       ),
      .wdata_i(wdata_i[bank]                     ),
      .be_i   (be_i[bank]                        ),
      .addr_i (addr_i[bank][$clog2(NumWords)-1:0])
    );
`else
  logic [NrBanks-1:0][8*StrbWidth-1:0] be_i_o;
  always_comb begin
    for(int i=0; i<StrbWidth; i++) begin
      be_i_o[bank][i*8 +: 8] = {8{be_i[bank][i]}};
    end
  end
 TS1N28HPCPUHDSVTB16X64M1SWBSO data_sram(
   .SLP  (1'b0),
   .SD   (1'b0),
   .CLK  (vrf_clk),
   .CEB  (!req_i[bank]),
   .WEB  (!wen_i[bank]),
   .CEBM (1'b1),
   .WEBM (1'b1),
   .A    (addr_i[bank][$clog2(NumWords)-1:0]),
   .D    (wdata_i[bank]),
   .BWEB (~be_i_o[bank]),
   .AM   ('0),
   .DM   ('0),
   .BWEBM('1),
   .BIST (1'b0),
   .RTSEL(2'b01),
   .WTSEL(2'b0),
   .Q    (rdata[bank]));
`endif
  end : gen_banks

  ///////////////////
  //  Multiplexer  //
  ///////////////////

  stream_xbar #(
    .NumInp   (NrBanks        ),
    .NumOut   (NrOperandQueues),
    .DataWidth(DataWidth      ),
    .AxiVldRdy('1             )
  ) i_vrf_mux (
    .clk_i  (clk_i          ),
    .rst_ni (rst_ni         ),
    .flush_i(1'b0           ),
    .rr_i   ('0             ),
    .data_i (rdata          ),
    .valid_i(rdata_valid_q  ),
    .ready_o(/* Unused */   ),
    .sel_i  (tgt_opqueue_q  ),
    .data_o (operand_o      ),
    .valid_o(operand_valid_o),
    .idx_o  (/* Unused */   ),
    .ready_i('1             ) // Always ready
  );

endmodule : vector_regfile
